library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity gameover_rom is
   Port (
       x_coord : in std_logic_vector(6 downto 0);
	   y_coord : in std_logic_vector(5 downto 0);
       rgb : out std_logic_vector(5 downto 0)
   );
end gameover_rom;


architecture Behavioral of gameover_rom is
signal total : std_logic_vector(12 downto 0);
begin
total <= y_coord & x_coord;
   process(total)
   begin
	case total is
       when "0001000010001" => rgb <= "000000";
        when "0001000010010" => rgb <= "000000";
        when "0001000010011" => rgb <= "000000";
        when "0001000010100" => rgb <= "000000";
        when "0001000011010" => rgb <= "000000";
        when "0001000011011" => rgb <= "000000";
        when "0001000011100" => rgb <= "000000";
        when "0001000011101" => rgb <= "000000";
        when "0001000011110" => rgb <= "000000";
        when "0001010001111" => rgb <= "000000";
        when "0001010010000" => rgb <= "000000";
        when "0001010010001" => rgb <= "100000";
        when "0001010010010" => rgb <= "100000";
        when "0001010010011" => rgb <= "100000";
        when "0001010010100" => rgb <= "100000";
        when "0001010010101" => rgb <= "000000";
        when "0001010010110" => rgb <= "000000";
        when "0001010011000" => rgb <= "000000";
        when "0001010011001" => rgb <= "000000";
        when "0001010011010" => rgb <= "101000";
        when "0001010011011" => rgb <= "101000";
        when "0001010011100" => rgb <= "101000";
        when "0001010011101" => rgb <= "101000";
        when "0001010011110" => rgb <= "101000";
        when "0001010011111" => rgb <= "000000";
        when "0001010100000" => rgb <= "000000";
        when "0001010100101" => rgb <= "000000";
        when "0001010100110" => rgb <= "000000";
        when "0001010100111" => rgb <= "000000";
        when "0001010110101" => rgb <= "000000";
        when "0001010110110" => rgb <= "000000";
        when "0001010110111" => rgb <= "000000";
        when "0001010111000" => rgb <= "000000";
        when "0001010111001" => rgb <= "000000";
        when "0001010111010" => rgb <= "000000";
        when "0001010111011" => rgb <= "000000";
        when "0001010111100" => rgb <= "000000";
        when "0001010111101" => rgb <= "000000";
        when "0001010111110" => rgb <= "000000";
        when "0001100001110" => rgb <= "000000";
        when "0001100001111" => rgb <= "100000";
        when "0001100010000" => rgb <= "100000";
        when "0001100010001" => rgb <= "100000";
        when "0001100010010" => rgb <= "100000";
        when "0001100010011" => rgb <= "100000";
        when "0001100010100" => rgb <= "100000";
        when "0001100010101" => rgb <= "100000";
        when "0001100010110" => rgb <= "000000";
        when "0001100010111" => rgb <= "000000";
        when "0001100011000" => rgb <= "101000";
        when "0001100011001" => rgb <= "101000";
        when "0001100011010" => rgb <= "101000";
        when "0001100011011" => rgb <= "101000";
        when "0001100011100" => rgb <= "101000";
        when "0001100011101" => rgb <= "101000";
        when "0001100011110" => rgb <= "101000";
        when "0001100011111" => rgb <= "101000";
        when "0001100100000" => rgb <= "101000";
        when "0001100100001" => rgb <= "000000";
        when "0001100100101" => rgb <= "000000";
        when "0001100100110" => rgb <= "001010";
        when "0001100100111" => rgb <= "001010";
        when "0001100101000" => rgb <= "000000";
        when "0001100101001" => rgb <= "000000";
        when "0001100110000" => rgb <= "000000";
        when "0001100110001" => rgb <= "000000";
        when "0001100110010" => rgb <= "000000";
        when "0001100110011" => rgb <= "000000";
        when "0001100110100" => rgb <= "000000";
        when "0001100110101" => rgb <= "100110";
        when "0001100110110" => rgb <= "100110";
        when "0001100110111" => rgb <= "100110";
        when "0001100111000" => rgb <= "100110";
        when "0001100111001" => rgb <= "100110";
        when "0001100111010" => rgb <= "100110";
        when "0001100111011" => rgb <= "100110";
        when "0001100111100" => rgb <= "100110";
        when "0001100111101" => rgb <= "100110";
        when "0001100111110" => rgb <= "000000";
        when "0001100111111" => rgb <= "000000";
        when "0001101000000" => rgb <= "000000";
        when "0001110001101" => rgb <= "000000";
        when "0001110001110" => rgb <= "100000";
        when "0001110001111" => rgb <= "100000";
        when "0001110010000" => rgb <= "100000";
        when "0001110010001" => rgb <= "100000";
        when "0001110010010" => rgb <= "100000";
        when "0001110010011" => rgb <= "100000";
        when "0001110010100" => rgb <= "100000";
        when "0001110010101" => rgb <= "100000";
        when "0001110010110" => rgb <= "100000";
        when "0001110010111" => rgb <= "000000";
        when "0001110011000" => rgb <= "101000";
        when "0001110011001" => rgb <= "101000";
        when "0001110011010" => rgb <= "101000";
        when "0001110011011" => rgb <= "101000";
        when "0001110011100" => rgb <= "101000";
        when "0001110011101" => rgb <= "101000";
        when "0001110011110" => rgb <= "101000";
        when "0001110011111" => rgb <= "101000";
        when "0001110100000" => rgb <= "101000";
        when "0001110100001" => rgb <= "101000";
        when "0001110100010" => rgb <= "000000";
        when "0001110100100" => rgb <= "000000";
        when "0001110100101" => rgb <= "001010";
        when "0001110100110" => rgb <= "001010";
        when "0001110100111" => rgb <= "001010";
        when "0001110101000" => rgb <= "001010";
        when "0001110101001" => rgb <= "000000";
        when "0001110101111" => rgb <= "000000";
        when "0001110110000" => rgb <= "001010";
        when "0001110110001" => rgb <= "001010";
        when "0001110110010" => rgb <= "000000";
        when "0001110110011" => rgb <= "000000";
        when "0001110110100" => rgb <= "100110";
        when "0001110110101" => rgb <= "100110";
        when "0001110110110" => rgb <= "100110";
        when "0001110110111" => rgb <= "100110";
        when "0001110111000" => rgb <= "100110";
        when "0001110111001" => rgb <= "100110";
        when "0001110111010" => rgb <= "100110";
        when "0001110111011" => rgb <= "100110";
        when "0001110111100" => rgb <= "100110";
        when "0001110111101" => rgb <= "100110";
        when "0001110111110" => rgb <= "100110";
        when "0001110111111" => rgb <= "100110";
        when "0001111000000" => rgb <= "000000";
        when "0001111000001" => rgb <= "000000";
        when "0010000001100" => rgb <= "000000";
        when "0010000001101" => rgb <= "000000";
        when "0010000001110" => rgb <= "100000";
        when "0010000001111" => rgb <= "100000";
        when "0010000010000" => rgb <= "100000";
        when "0010000010001" => rgb <= "100000";
        when "0010000010010" => rgb <= "000000";
        when "0010000010011" => rgb <= "000000";
        when "0010000010100" => rgb <= "100000";
        when "0010000010101" => rgb <= "100000";
        when "0010000010110" => rgb <= "100000";
        when "0010000010111" => rgb <= "000000";
        when "0010000011000" => rgb <= "101000";
        when "0010000011001" => rgb <= "101000";
        when "0010000011010" => rgb <= "101000";
        when "0010000011011" => rgb <= "101000";
        when "0010000011100" => rgb <= "101000";
        when "0010000011101" => rgb <= "101000";
        when "0010000011110" => rgb <= "101000";
        when "0010000011111" => rgb <= "101000";
        when "0010000100000" => rgb <= "101000";
        when "0010000100001" => rgb <= "101000";
        when "0010000100010" => rgb <= "000000";
        when "0010000100011" => rgb <= "000000";
        when "0010000100100" => rgb <= "000000";
        when "0010000100101" => rgb <= "001010";
        when "0010000100110" => rgb <= "001010";
        when "0010000100111" => rgb <= "001010";
        when "0010000101000" => rgb <= "001010";
        when "0010000101001" => rgb <= "001010";
        when "0010000101010" => rgb <= "000000";
        when "0010000101110" => rgb <= "000000";
        when "0010000101111" => rgb <= "001010";
        when "0010000110000" => rgb <= "001010";
        when "0010000110001" => rgb <= "001010";
        when "0010000110010" => rgb <= "001010";
        when "0010000110011" => rgb <= "000000";
        when "0010000110100" => rgb <= "100110";
        when "0010000110101" => rgb <= "100110";
        when "0010000110110" => rgb <= "100110";
        when "0010000110111" => rgb <= "100110";
        when "0010000111000" => rgb <= "100110";
        when "0010000111001" => rgb <= "100110";
        when "0010000111010" => rgb <= "100110";
        when "0010000111011" => rgb <= "100110";
        when "0010000111100" => rgb <= "100110";
        when "0010000111101" => rgb <= "100110";
        when "0010000111110" => rgb <= "100110";
        when "0010000111111" => rgb <= "100110";
        when "0010001000000" => rgb <= "100110";
        when "0010001000001" => rgb <= "000000";
        when "0010010001100" => rgb <= "000000";
        when "0010010001101" => rgb <= "100000";
        when "0010010001110" => rgb <= "100000";
        when "0010010001111" => rgb <= "100000";
        when "0010010010000" => rgb <= "100000";
        when "0010010010001" => rgb <= "000000";
        when "0010010010100" => rgb <= "000000";
        when "0010010010101" => rgb <= "100000";
        when "0010010010110" => rgb <= "100000";
        when "0010010010111" => rgb <= "000000";
        when "0010010011000" => rgb <= "101000";
        when "0010010011001" => rgb <= "000000";
        when "0010010011010" => rgb <= "000000";
        when "0010010011011" => rgb <= "000000";
        when "0010010011100" => rgb <= "000000";
        when "0010010011101" => rgb <= "101000";
        when "0010010011110" => rgb <= "000000";
        when "0010010011111" => rgb <= "000000";
        when "0010010100000" => rgb <= "000000";
        when "0010010100001" => rgb <= "000000";
        when "0010010100010" => rgb <= "101000";
        when "0010010100011" => rgb <= "000000";
        when "0010010100100" => rgb <= "000000";
        when "0010010100101" => rgb <= "001010";
        when "0010010100110" => rgb <= "001010";
        when "0010010100111" => rgb <= "001010";
        when "0010010101000" => rgb <= "001010";
        when "0010010101001" => rgb <= "001010";
        when "0010010101010" => rgb <= "000000";
        when "0010010101011" => rgb <= "000000";
        when "0010010101101" => rgb <= "000000";
        when "0010010101110" => rgb <= "001010";
        when "0010010101111" => rgb <= "001010";
        when "0010010110000" => rgb <= "001010";
        when "0010010110001" => rgb <= "001010";
        when "0010010110010" => rgb <= "001010";
        when "0010010110011" => rgb <= "000000";
        when "0010010110100" => rgb <= "000000";
        when "0010010110101" => rgb <= "100110";
        when "0010010110110" => rgb <= "100110";
        when "0010010110111" => rgb <= "100110";
        when "0010010111000" => rgb <= "100110";
        when "0010010111001" => rgb <= "000000";
        when "0010010111010" => rgb <= "000000";
        when "0010010111011" => rgb <= "000000";
        when "0010010111100" => rgb <= "000000";
        when "0010010111101" => rgb <= "000000";
        when "0010010111110" => rgb <= "000000";
        when "0010010111111" => rgb <= "000000";
        when "0010011000000" => rgb <= "000000";
        when "0010011000001" => rgb <= "000000";
        when "0010100001011" => rgb <= "000000";
        when "0010100001100" => rgb <= "000000";
        when "0010100001101" => rgb <= "100000";
        when "0010100001110" => rgb <= "100000";
        when "0010100001111" => rgb <= "100000";
        when "0010100010000" => rgb <= "100000";
        when "0010100010001" => rgb <= "000000";
        when "0010100010101" => rgb <= "000000";
        when "0010100010110" => rgb <= "000000";
        when "0010100010111" => rgb <= "101000";
        when "0010100011000" => rgb <= "101000";
        when "0010100011001" => rgb <= "000000";
        when "0010100011010" => rgb <= "000000";
        when "0010100011011" => rgb <= "101010";
        when "0010100011100" => rgb <= "000000";
        when "0010100011101" => rgb <= "101000";
        when "0010100011110" => rgb <= "000000";
        when "0010100011111" => rgb <= "000000";
        when "0010100100000" => rgb <= "101010";
        when "0010100100001" => rgb <= "000000";
        when "0010100100010" => rgb <= "101000";
        when "0010100100011" => rgb <= "101000";
        when "0010100100100" => rgb <= "000000";
        when "0010100100101" => rgb <= "001010";
        when "0010100100110" => rgb <= "001010";
        when "0010100100111" => rgb <= "001010";
        when "0010100101000" => rgb <= "001010";
        when "0010100101001" => rgb <= "001010";
        when "0010100101010" => rgb <= "001010";
        when "0010100101011" => rgb <= "000000";
        when "0010100101101" => rgb <= "000000";
        when "0010100101110" => rgb <= "001010";
        when "0010100101111" => rgb <= "001010";
        when "0010100110000" => rgb <= "001010";
        when "0010100110001" => rgb <= "001010";
        when "0010100110010" => rgb <= "001010";
        when "0010100110011" => rgb <= "001010";
        when "0010100110100" => rgb <= "000000";
        when "0010100110101" => rgb <= "100110";
        when "0010100110110" => rgb <= "100110";
        when "0010100110111" => rgb <= "100110";
        when "0010100111000" => rgb <= "100110";
        when "0010100111001" => rgb <= "000000";
        when "0010110001011" => rgb <= "000000";
        when "0010110001100" => rgb <= "100000";
        when "0010110001101" => rgb <= "100000";
        when "0010110001110" => rgb <= "100000";
        when "0010110001111" => rgb <= "100000";
        when "0010110010000" => rgb <= "000000";
        when "0010110010110" => rgb <= "000000";
        when "0010110010111" => rgb <= "101000";
        when "0010110011000" => rgb <= "101000";
        when "0010110011001" => rgb <= "000000";
        when "0010110011010" => rgb <= "101010";
        when "0010110011011" => rgb <= "101010";
        when "0010110011100" => rgb <= "000000";
        when "0010110011101" => rgb <= "101000";
        when "0010110011110" => rgb <= "000000";
        when "0010110011111" => rgb <= "101010";
        when "0010110100000" => rgb <= "101010";
        when "0010110100001" => rgb <= "000000";
        when "0010110100010" => rgb <= "101000";
        when "0010110100011" => rgb <= "101000";
        when "0010110100100" => rgb <= "000000";
        when "0010110100101" => rgb <= "001010";
        when "0010110100110" => rgb <= "001010";
        when "0010110100111" => rgb <= "001010";
        when "0010110101000" => rgb <= "001010";
        when "0010110101001" => rgb <= "001010";
        when "0010110101010" => rgb <= "001010";
        when "0010110101011" => rgb <= "001010";
        when "0010110101100" => rgb <= "000000";
        when "0010110101101" => rgb <= "000000";
        when "0010110101110" => rgb <= "001010";
        when "0010110101111" => rgb <= "001010";
        when "0010110110000" => rgb <= "001010";
        when "0010110110001" => rgb <= "001010";
        when "0010110110010" => rgb <= "001010";
        when "0010110110011" => rgb <= "001010";
        when "0010110110100" => rgb <= "000000";
        when "0010110110101" => rgb <= "100110";
        when "0010110110110" => rgb <= "100110";
        when "0010110110111" => rgb <= "100110";
        when "0010110111000" => rgb <= "100110";
        when "0010110111001" => rgb <= "000000";
        when "0010110111010" => rgb <= "000000";
        when "0010110111011" => rgb <= "000000";
        when "0011000001011" => rgb <= "000000";
        when "0011000001100" => rgb <= "100000";
        when "0011000001101" => rgb <= "100000";
        when "0011000001110" => rgb <= "100000";
        when "0011000001111" => rgb <= "100000";
        when "0011000010000" => rgb <= "000000";
        when "0011000010110" => rgb <= "000000";
        when "0011000010111" => rgb <= "101000";
        when "0011000011000" => rgb <= "101000";
        when "0011000011001" => rgb <= "000000";
        when "0011000011010" => rgb <= "000000";
        when "0011000011011" => rgb <= "000000";
        when "0011000011100" => rgb <= "000000";
        when "0011000011101" => rgb <= "101000";
        when "0011000011110" => rgb <= "000000";
        when "0011000011111" => rgb <= "000000";
        when "0011000100000" => rgb <= "000000";
        when "0011000100001" => rgb <= "000000";
        when "0011000100010" => rgb <= "101000";
        when "0011000100011" => rgb <= "101000";
        when "0011000100100" => rgb <= "000000";
        when "0011000100101" => rgb <= "001010";
        when "0011000100110" => rgb <= "001010";
        when "0011000100111" => rgb <= "001010";
        when "0011000101000" => rgb <= "001010";
        when "0011000101001" => rgb <= "001010";
        when "0011000101010" => rgb <= "001010";
        when "0011000101011" => rgb <= "001010";
        when "0011000101100" => rgb <= "001010";
        when "0011000101101" => rgb <= "001010";
        when "0011000101110" => rgb <= "001010";
        when "0011000101111" => rgb <= "001010";
        when "0011000110000" => rgb <= "001010";
        when "0011000110001" => rgb <= "001010";
        when "0011000110010" => rgb <= "001010";
        when "0011000110011" => rgb <= "001010";
        when "0011000110100" => rgb <= "000000";
        when "0011000110101" => rgb <= "100110";
        when "0011000110110" => rgb <= "100110";
        when "0011000110111" => rgb <= "100110";
        when "0011000111000" => rgb <= "100110";
        when "0011000111001" => rgb <= "100110";
        when "0011000111010" => rgb <= "100110";
        when "0011000111011" => rgb <= "100110";
        when "0011000111100" => rgb <= "000000";
        when "0011000111101" => rgb <= "000000";
        when "0011010001011" => rgb <= "000000";
        when "0011010001100" => rgb <= "100000";
        when "0011010001101" => rgb <= "100000";
        when "0011010001110" => rgb <= "100000";
        when "0011010001111" => rgb <= "100000";
        when "0011010010000" => rgb <= "000000";
        when "0011010010110" => rgb <= "000000";
        when "0011010010111" => rgb <= "101000";
        when "0011010011000" => rgb <= "101000";
        when "0011010011001" => rgb <= "101000";
        when "0011010011010" => rgb <= "101000";
        when "0011010011011" => rgb <= "101000";
        when "0011010011100" => rgb <= "101000";
        when "0011010011101" => rgb <= "101000";
        when "0011010011110" => rgb <= "101000";
        when "0011010011111" => rgb <= "101000";
        when "0011010100000" => rgb <= "101000";
        when "0011010100001" => rgb <= "101000";
        when "0011010100010" => rgb <= "101000";
        when "0011010100011" => rgb <= "101000";
        when "0011010100100" => rgb <= "101000";
        when "0011010100101" => rgb <= "000000";
        when "0011010100110" => rgb <= "001010";
        when "0011010100111" => rgb <= "001010";
        when "0011010101000" => rgb <= "001010";
        when "0011010101001" => rgb <= "001010";
        when "0011010101010" => rgb <= "001010";
        when "0011010101011" => rgb <= "001010";
        when "0011010101100" => rgb <= "001010";
        when "0011010101101" => rgb <= "001010";
        when "0011010101110" => rgb <= "001010";
        when "0011010101111" => rgb <= "001010";
        when "0011010110000" => rgb <= "001010";
        when "0011010110001" => rgb <= "001010";
        when "0011010110010" => rgb <= "001010";
        when "0011010110011" => rgb <= "001010";
        when "0011010110100" => rgb <= "000000";
        when "0011010110101" => rgb <= "100110";
        when "0011010110110" => rgb <= "100110";
        when "0011010110111" => rgb <= "100110";
        when "0011010111000" => rgb <= "100110";
        when "0011010111001" => rgb <= "100110";
        when "0011010111010" => rgb <= "100110";
        when "0011010111011" => rgb <= "100110";
        when "0011010111100" => rgb <= "100110";
        when "0011010111101" => rgb <= "000000";
        when "0011100001100" => rgb <= "000000";
        when "0011100001101" => rgb <= "100000";
        when "0011100001110" => rgb <= "100000";
        when "0011100001111" => rgb <= "100000";
        when "0011100010000" => rgb <= "000000";
        when "0011100010101" => rgb <= "000000";
        when "0011100010110" => rgb <= "000000";
        when "0011100010111" => rgb <= "000000";
        when "0011100011000" => rgb <= "101000";
        when "0011100011001" => rgb <= "101000";
        when "0011100011010" => rgb <= "101000";
        when "0011100011011" => rgb <= "101000";
        when "0011100011100" => rgb <= "101000";
        when "0011100011101" => rgb <= "101000";
        when "0011100011110" => rgb <= "101000";
        when "0011100011111" => rgb <= "101000";
        when "0011100100000" => rgb <= "101000";
        when "0011100100001" => rgb <= "101000";
        when "0011100100010" => rgb <= "101000";
        when "0011100100011" => rgb <= "101000";
        when "0011100100100" => rgb <= "101000";
        when "0011100100101" => rgb <= "000000";
        when "0011100100110" => rgb <= "001010";
        when "0011100100111" => rgb <= "001010";
        when "0011100101000" => rgb <= "001010";
        when "0011100101001" => rgb <= "001010";
        when "0011100101010" => rgb <= "000000";
        when "0011100101011" => rgb <= "001010";
        when "0011100101100" => rgb <= "001010";
        when "0011100101101" => rgb <= "001010";
        when "0011100101110" => rgb <= "001010";
        when "0011100101111" => rgb <= "000000";
        when "0011100110000" => rgb <= "001010";
        when "0011100110001" => rgb <= "001010";
        when "0011100110010" => rgb <= "001010";
        when "0011100110011" => rgb <= "001010";
        when "0011100110100" => rgb <= "001010";
        when "0011100110101" => rgb <= "000000";
        when "0011100110110" => rgb <= "100110";
        when "0011100110111" => rgb <= "100110";
        when "0011100111000" => rgb <= "100110";
        when "0011100111001" => rgb <= "100110";
        when "0011100111010" => rgb <= "000000";
        when "0011100111011" => rgb <= "000000";
        when "0011100111100" => rgb <= "000000";
        when "0011100111101" => rgb <= "000000";
        when "0011110001100" => rgb <= "000000";
        when "0011110001101" => rgb <= "100000";
        when "0011110001110" => rgb <= "100000";
        when "0011110001111" => rgb <= "100000";
        when "0011110010000" => rgb <= "000000";
        when "0011110010011" => rgb <= "000000";
        when "0011110010100" => rgb <= "000000";
        when "0011110010101" => rgb <= "100000";
        when "0011110010110" => rgb <= "100000";
        when "0011110010111" => rgb <= "000000";
        when "0011110011000" => rgb <= "000000";
        when "0011110011001" => rgb <= "101000";
        when "0011110011010" => rgb <= "101000";
        when "0011110011011" => rgb <= "101000";
        when "0011110011100" => rgb <= "101000";
        when "0011110011101" => rgb <= "101000";
        when "0011110011110" => rgb <= "101000";
        when "0011110011111" => rgb <= "101000";
        when "0011110100000" => rgb <= "101000";
        when "0011110100001" => rgb <= "101000";
        when "0011110100010" => rgb <= "101000";
        when "0011110100011" => rgb <= "101000";
        when "0011110100100" => rgb <= "101000";
        when "0011110100101" => rgb <= "000000";
        when "0011110100110" => rgb <= "001010";
        when "0011110100111" => rgb <= "001010";
        when "0011110101000" => rgb <= "001010";
        when "0011110101001" => rgb <= "000000";
        when "0011110101010" => rgb <= "000000";
        when "0011110101011" => rgb <= "001010";
        when "0011110101100" => rgb <= "001010";
        when "0011110101101" => rgb <= "001010";
        when "0011110101110" => rgb <= "000000";
        when "0011110110000" => rgb <= "000000";
        when "0011110110001" => rgb <= "001010";
        when "0011110110010" => rgb <= "001010";
        when "0011110110011" => rgb <= "001010";
        when "0011110110100" => rgb <= "001010";
        when "0011110110101" => rgb <= "000000";
        when "0011110110110" => rgb <= "100110";
        when "0011110110111" => rgb <= "100110";
        when "0011110111000" => rgb <= "100110";
        when "0011110111001" => rgb <= "100110";
        when "0011110111010" => rgb <= "000000";
        when "0100000001100" => rgb <= "000000";
        when "0100000001101" => rgb <= "100000";
        when "0100000001110" => rgb <= "100000";
        when "0100000001111" => rgb <= "100000";
        when "0100000010000" => rgb <= "000000";
        when "0100000010011" => rgb <= "000000";
        when "0100000010100" => rgb <= "100000";
        when "0100000010101" => rgb <= "100000";
        when "0100000010110" => rgb <= "100000";
        when "0100000010111" => rgb <= "100000";
        when "0100000011000" => rgb <= "100000";
        when "0100000011001" => rgb <= "000000";
        when "0100000011010" => rgb <= "101000";
        when "0100000011011" => rgb <= "101000";
        when "0100000011100" => rgb <= "101000";
        when "0100000011101" => rgb <= "101000";
        when "0100000011110" => rgb <= "101000";
        when "0100000011111" => rgb <= "101000";
        when "0100000100000" => rgb <= "101000";
        when "0100000100001" => rgb <= "101000";
        when "0100000100010" => rgb <= "101000";
        when "0100000100011" => rgb <= "101000";
        when "0100000100100" => rgb <= "101000";
        when "0100000100101" => rgb <= "000000";
        when "0100000100110" => rgb <= "001010";
        when "0100000100111" => rgb <= "001010";
        when "0100000101000" => rgb <= "001010";
        when "0100000101001" => rgb <= "000000";
        when "0100000101010" => rgb <= "000000";
        when "0100000101011" => rgb <= "000000";
        when "0100000101100" => rgb <= "000000";
        when "0100000101101" => rgb <= "000000";
        when "0100000101110" => rgb <= "000000";
        when "0100000110000" => rgb <= "000000";
        when "0100000110001" => rgb <= "001010";
        when "0100000110010" => rgb <= "001010";
        when "0100000110011" => rgb <= "001010";
        when "0100000110100" => rgb <= "001010";
        when "0100000110101" => rgb <= "000000";
        when "0100000110110" => rgb <= "100110";
        when "0100000110111" => rgb <= "100110";
        when "0100000111000" => rgb <= "100110";
        when "0100000111001" => rgb <= "100110";
        when "0100000111010" => rgb <= "000000";
        when "0100010001101" => rgb <= "000000";
        when "0100010001110" => rgb <= "100000";
        when "0100010001111" => rgb <= "100000";
        when "0100010010000" => rgb <= "100000";
        when "0100010010001" => rgb <= "000000";
        when "0100010010100" => rgb <= "000000";
        when "0100010010101" => rgb <= "000000";
        when "0100010010110" => rgb <= "000000";
        when "0100010010111" => rgb <= "100000";
        when "0100010011000" => rgb <= "100000";
        when "0100010011001" => rgb <= "000000";
        when "0100010011010" => rgb <= "101000";
        when "0100010011011" => rgb <= "101000";
        when "0100010011100" => rgb <= "101000";
        when "0100010011101" => rgb <= "101000";
        when "0100010011110" => rgb <= "101000";
        when "0100010011111" => rgb <= "101000";
        when "0100010100000" => rgb <= "101000";
        when "0100010100001" => rgb <= "101000";
        when "0100010100010" => rgb <= "101000";
        when "0100010100011" => rgb <= "101000";
        when "0100010100100" => rgb <= "101000";
        when "0100010100101" => rgb <= "000000";
        when "0100010100110" => rgb <= "001010";
        when "0100010100111" => rgb <= "001010";
        when "0100010101000" => rgb <= "001010";
        when "0100010101001" => rgb <= "000000";
        when "0100010110000" => rgb <= "000000";
        when "0100010110001" => rgb <= "001010";
        when "0100010110010" => rgb <= "001010";
        when "0100010110011" => rgb <= "001010";
        when "0100010110100" => rgb <= "001010";
        when "0100010110101" => rgb <= "000000";
        when "0100010110110" => rgb <= "100110";
        when "0100010110111" => rgb <= "100110";
        when "0100010111000" => rgb <= "100110";
        when "0100010111001" => rgb <= "100110";
        when "0100010111010" => rgb <= "000000";
        when "0100010111011" => rgb <= "000000";
        when "0100010111100" => rgb <= "000000";
        when "0100010111101" => rgb <= "000000";
        when "0100010111110" => rgb <= "000000";
        when "0100010111111" => rgb <= "000000";
        when "0100011000000" => rgb <= "000000";
        when "0100011000001" => rgb <= "000000";
        when "0100011000010" => rgb <= "000000";
        when "0100100001101" => rgb <= "000000";
        when "0100100001110" => rgb <= "100000";
        when "0100100001111" => rgb <= "100000";
        when "0100100010000" => rgb <= "100000";
        when "0100100010001" => rgb <= "100000";
        when "0100100010010" => rgb <= "000000";
        when "0100100010011" => rgb <= "000000";
        when "0100100010101" => rgb <= "000000";
        when "0100100010110" => rgb <= "100000";
        when "0100100010111" => rgb <= "100000";
        when "0100100011000" => rgb <= "100000";
        when "0100100011001" => rgb <= "000000";
        when "0100100011010" => rgb <= "101000";
        when "0100100011011" => rgb <= "101000";
        when "0100100011100" => rgb <= "101000";
        when "0100100011101" => rgb <= "101000";
        when "0100100011110" => rgb <= "101000";
        when "0100100011111" => rgb <= "101000";
        when "0100100100000" => rgb <= "101000";
        when "0100100100001" => rgb <= "101000";
        when "0100100100010" => rgb <= "101000";
        when "0100100100011" => rgb <= "101000";
        when "0100100100100" => rgb <= "101000";
        when "0100100100101" => rgb <= "000000";
        when "0100100100110" => rgb <= "001010";
        when "0100100100111" => rgb <= "001010";
        when "0100100101000" => rgb <= "001010";
        when "0100100101001" => rgb <= "000000";
        when "0100100110000" => rgb <= "000000";
        when "0100100110001" => rgb <= "001010";
        when "0100100110010" => rgb <= "001010";
        when "0100100110011" => rgb <= "001010";
        when "0100100110100" => rgb <= "001010";
        when "0100100110101" => rgb <= "000000";
        when "0100100110110" => rgb <= "100110";
        when "0100100110111" => rgb <= "100110";
        when "0100100111000" => rgb <= "100110";
        when "0100100111001" => rgb <= "100110";
        when "0100100111010" => rgb <= "100110";
        when "0100100111011" => rgb <= "100110";
        when "0100100111100" => rgb <= "100110";
        when "0100100111101" => rgb <= "100110";
        when "0100100111110" => rgb <= "100110";
        when "0100100111111" => rgb <= "100110";
        when "0100101000000" => rgb <= "100110";
        when "0100101000001" => rgb <= "100110";
        when "0100101000010" => rgb <= "000000";
        when "0100110001110" => rgb <= "000000";
        when "0100110001111" => rgb <= "100000";
        when "0100110010000" => rgb <= "100000";
        when "0100110010001" => rgb <= "100000";
        when "0100110010010" => rgb <= "100000";
        when "0100110010011" => rgb <= "100000";
        when "0100110010100" => rgb <= "000000";
        when "0100110010101" => rgb <= "000000";
        when "0100110010110" => rgb <= "100000";
        when "0100110010111" => rgb <= "100000";
        when "0100110011000" => rgb <= "100000";
        when "0100110011001" => rgb <= "000000";
        when "0100110011010" => rgb <= "101000";
        when "0100110011011" => rgb <= "101000";
        when "0100110011100" => rgb <= "101000";
        when "0100110011101" => rgb <= "101000";
        when "0100110011110" => rgb <= "000000";
        when "0100110011111" => rgb <= "101000";
        when "0100110100000" => rgb <= "101000";
        when "0100110100001" => rgb <= "101000";
        when "0100110100010" => rgb <= "101000";
        when "0100110100011" => rgb <= "101000";
        when "0100110100100" => rgb <= "101000";
        when "0100110100101" => rgb <= "000000";
        when "0100110100110" => rgb <= "001010";
        when "0100110100111" => rgb <= "001010";
        when "0100110101000" => rgb <= "001010";
        when "0100110101001" => rgb <= "000000";
        when "0100110110000" => rgb <= "000000";
        when "0100110110001" => rgb <= "001010";
        when "0100110110010" => rgb <= "001010";
        when "0100110110011" => rgb <= "001010";
        when "0100110110100" => rgb <= "001010";
        when "0100110110101" => rgb <= "000000";
        when "0100110110110" => rgb <= "100110";
        when "0100110110111" => rgb <= "100110";
        when "0100110111000" => rgb <= "100110";
        when "0100110111001" => rgb <= "100110";
        when "0100110111010" => rgb <= "100110";
        when "0100110111011" => rgb <= "100110";
        when "0100110111100" => rgb <= "100110";
        when "0100110111101" => rgb <= "100110";
        when "0100110111110" => rgb <= "100110";
        when "0100110111111" => rgb <= "100110";
        when "0100111000000" => rgb <= "100110";
        when "0100111000001" => rgb <= "100110";
        when "0100111000010" => rgb <= "000000";
        when "0101000001110" => rgb <= "000000";
        when "0101000001111" => rgb <= "000000";
        when "0101000010000" => rgb <= "100000";
        when "0101000010001" => rgb <= "100000";
        when "0101000010010" => rgb <= "100000";
        when "0101000010011" => rgb <= "100000";
        when "0101000010100" => rgb <= "100000";
        when "0101000010101" => rgb <= "100000";
        when "0101000010110" => rgb <= "100000";
        when "0101000010111" => rgb <= "100000";
        when "0101000011000" => rgb <= "000000";
        when "0101000011001" => rgb <= "000000";
        when "0101000011010" => rgb <= "101000";
        when "0101000011011" => rgb <= "000000";
        when "0101000011100" => rgb <= "101000";
        when "0101000011101" => rgb <= "101000";
        when "0101000011110" => rgb <= "000000";
        when "0101000011111" => rgb <= "000000";
        when "0101000100000" => rgb <= "101000";
        when "0101000100001" => rgb <= "101000";
        when "0101000100010" => rgb <= "000000";
        when "0101000100011" => rgb <= "101000";
        when "0101000100100" => rgb <= "101000";
        when "0101000100101" => rgb <= "000000";
        when "0101000100110" => rgb <= "001010";
        when "0101000100111" => rgb <= "001010";
        when "0101000101000" => rgb <= "000000";
        when "0101000101001" => rgb <= "000000";
        when "0101000110000" => rgb <= "000000";
        when "0101000110001" => rgb <= "000000";
        when "0101000110010" => rgb <= "001010";
        when "0101000110011" => rgb <= "001010";
        when "0101000110100" => rgb <= "001010";
        when "0101000110101" => rgb <= "000000";
        when "0101000110110" => rgb <= "100110";
        when "0101000110111" => rgb <= "100110";
        when "0101000111000" => rgb <= "100110";
        when "0101000111001" => rgb <= "100110";
        when "0101000111010" => rgb <= "100110";
        when "0101000111011" => rgb <= "100110";
        when "0101000111100" => rgb <= "100110";
        when "0101000111101" => rgb <= "100110";
        when "0101000111110" => rgb <= "100110";
        when "0101000111111" => rgb <= "100110";
        when "0101001000000" => rgb <= "100110";
        when "0101001000001" => rgb <= "000000";
        when "0101001000010" => rgb <= "000000";
        when "0101010001111" => rgb <= "000000";
        when "0101010010000" => rgb <= "000000";
        when "0101010010001" => rgb <= "100000";
        when "0101010010010" => rgb <= "100000";
        when "0101010010011" => rgb <= "100000";
        when "0101010010100" => rgb <= "100000";
        when "0101010010101" => rgb <= "100000";
        when "0101010010110" => rgb <= "100000";
        when "0101010010111" => rgb <= "000000";
        when "0101010011001" => rgb <= "000000";
        when "0101010011010" => rgb <= "000000";
        when "0101010011011" => rgb <= "000000";
        when "0101010011100" => rgb <= "101000";
        when "0101010011101" => rgb <= "000000";
        when "0101010011110" => rgb <= "000000";
        when "0101010011111" => rgb <= "000000";
        when "0101010100000" => rgb <= "000000";
        when "0101010100001" => rgb <= "101000";
        when "0101010100010" => rgb <= "000000";
        when "0101010100011" => rgb <= "000000";
        when "0101010100100" => rgb <= "101000";
        when "0101010100101" => rgb <= "000000";
        when "0101010100110" => rgb <= "000000";
        when "0101010100111" => rgb <= "000000";
        when "0101010101000" => rgb <= "000000";
        when "0101010110001" => rgb <= "000000";
        when "0101010110010" => rgb <= "000000";
        when "0101010110011" => rgb <= "000000";
        when "0101010110100" => rgb <= "000000";
        when "0101010110101" => rgb <= "000000";
        when "0101010110110" => rgb <= "000000";
        when "0101010110111" => rgb <= "000000";
        when "0101010111000" => rgb <= "000000";
        when "0101010111001" => rgb <= "000000";
        when "0101010111010" => rgb <= "000000";
        when "0101010111011" => rgb <= "000000";
        when "0101010111100" => rgb <= "000000";
        when "0101010111101" => rgb <= "000000";
        when "0101010111110" => rgb <= "000000";
        when "0101010111111" => rgb <= "000000";
        when "0101011000000" => rgb <= "000000";
        when "0101011000001" => rgb <= "000000";
        when "0101100010001" => rgb <= "000000";
        when "0101100010010" => rgb <= "000000";
        when "0101100010011" => rgb <= "000000";
        when "0101100010100" => rgb <= "000000";
        when "0101100010101" => rgb <= "000000";
        when "0101100010110" => rgb <= "000000";
        when "0101100011010" => rgb <= "000000";
        when "0101100011100" => rgb <= "000000";
        when "0101100011101" => rgb <= "000000";
        when "0101100100001" => rgb <= "000000";
        when "0101100100100" => rgb <= "000000";
        when "0110010010011" => rgb <= "000000";
        when "0110010010100" => rgb <= "000000";
        when "0110010010101" => rgb <= "000000";
        when "0110010010110" => rgb <= "000000";
        when "0110010011010" => rgb <= "000000";
        when "0110010011011" => rgb <= "000000";
        when "0110010011100" => rgb <= "000000";
        when "0110010101001" => rgb <= "000000";
        when "0110100010001" => rgb <= "000000";
        when "0110100010010" => rgb <= "000000";
        when "0110100010011" => rgb <= "101000";
        when "0110100010100" => rgb <= "101000";
        when "0110100010101" => rgb <= "101000";
        when "0110100010110" => rgb <= "101000";
        when "0110100010111" => rgb <= "000000";
        when "0110100011000" => rgb <= "000000";
        when "0110100011001" => rgb <= "000000";
        when "0110100011010" => rgb <= "000000";
        when "0110100011011" => rgb <= "100110";
        when "0110100011100" => rgb <= "100110";
        when "0110100011101" => rgb <= "000000";
        when "0110100011110" => rgb <= "000000";
        when "0110100100111" => rgb <= "000000";
        when "0110100101000" => rgb <= "000000";
        when "0110100101001" => rgb <= "100110";
        when "0110100101010" => rgb <= "000000";
        when "0110100110110" => rgb <= "000000";
        when "0110100110111" => rgb <= "000000";
        when "0110100111000" => rgb <= "000000";
        when "0110100111001" => rgb <= "000000";
        when "0110100111010" => rgb <= "000000";
        when "0110100111011" => rgb <= "000000";
        when "0110100111100" => rgb <= "000000";
        when "0110100111101" => rgb <= "000000";
        when "0110110001111" => rgb <= "000000";
        when "0110110010000" => rgb <= "000000";
        when "0110110010001" => rgb <= "101000";
        when "0110110010010" => rgb <= "101000";
        when "0110110010011" => rgb <= "101000";
        when "0110110010100" => rgb <= "101000";
        when "0110110010101" => rgb <= "101000";
        when "0110110010110" => rgb <= "101000";
        when "0110110010111" => rgb <= "101000";
        when "0110110011000" => rgb <= "101000";
        when "0110110011001" => rgb <= "101000";
        when "0110110011010" => rgb <= "000000";
        when "0110110011011" => rgb <= "100110";
        when "0110110011100" => rgb <= "100110";
        when "0110110011101" => rgb <= "100110";
        when "0110110011110" => rgb <= "000000";
        when "0110110011111" => rgb <= "000000";
        when "0110110100110" => rgb <= "000000";
        when "0110110100111" => rgb <= "000000";
        when "0110110101000" => rgb <= "100110";
        when "0110110101001" => rgb <= "100110";
        when "0110110101010" => rgb <= "100110";
        when "0110110101011" => rgb <= "000000";
        when "0110110101100" => rgb <= "000000";
        when "0110110101101" => rgb <= "000000";
        when "0110110101110" => rgb <= "000000";
        when "0110110101111" => rgb <= "000000";
        when "0110110110000" => rgb <= "000000";
        when "0110110110001" => rgb <= "000000";
        when "0110110110010" => rgb <= "000000";
        when "0110110110101" => rgb <= "000000";
        when "0110110110110" => rgb <= "101000";
        when "0110110110111" => rgb <= "101000";
        when "0110110111000" => rgb <= "101000";
        when "0110110111001" => rgb <= "101000";
        when "0110110111010" => rgb <= "101000";
        when "0110110111011" => rgb <= "101000";
        when "0110110111100" => rgb <= "101000";
        when "0110110111101" => rgb <= "101000";
        when "0110110111110" => rgb <= "000000";
        when "0110110111111" => rgb <= "000000";
        when "0111000001110" => rgb <= "000000";
        when "0111000001111" => rgb <= "000000";
        when "0111000010000" => rgb <= "101000";
        when "0111000010001" => rgb <= "101000";
        when "0111000010010" => rgb <= "101000";
        when "0111000010011" => rgb <= "101000";
        when "0111000010100" => rgb <= "101000";
        when "0111000010101" => rgb <= "101000";
        when "0111000010110" => rgb <= "101000";
        when "0111000010111" => rgb <= "101000";
        when "0111000011000" => rgb <= "101000";
        when "0111000011001" => rgb <= "101000";
        when "0111000011010" => rgb <= "000000";
        when "0111000011011" => rgb <= "100110";
        when "0111000011100" => rgb <= "100110";
        when "0111000011101" => rgb <= "100110";
        when "0111000011110" => rgb <= "100110";
        when "0111000011111" => rgb <= "000000";
        when "0111000100110" => rgb <= "000000";
        when "0111000100111" => rgb <= "100110";
        when "0111000101000" => rgb <= "100110";
        when "0111000101001" => rgb <= "100110";
        when "0111000101010" => rgb <= "000000";
        when "0111000101011" => rgb <= "000000";
        when "0111000101100" => rgb <= "100000";
        when "0111000101101" => rgb <= "100000";
        when "0111000101110" => rgb <= "100000";
        when "0111000101111" => rgb <= "100000";
        when "0111000110000" => rgb <= "100000";
        when "0111000110001" => rgb <= "100000";
        when "0111000110010" => rgb <= "100000";
        when "0111000110011" => rgb <= "000000";
        when "0111000110100" => rgb <= "000000";
        when "0111000110101" => rgb <= "000000";
        when "0111000110110" => rgb <= "101000";
        when "0111000110111" => rgb <= "101000";
        when "0111000111000" => rgb <= "101000";
        when "0111000111001" => rgb <= "101000";
        when "0111000111010" => rgb <= "101000";
        when "0111000111011" => rgb <= "101000";
        when "0111000111100" => rgb <= "101000";
        when "0111000111101" => rgb <= "101000";
        when "0111000111110" => rgb <= "101000";
        when "0111000111111" => rgb <= "000000";
        when "0111001000000" => rgb <= "000000";
        when "0111010001110" => rgb <= "000000";
        when "0111010001111" => rgb <= "101000";
        when "0111010010000" => rgb <= "101000";
        when "0111010010001" => rgb <= "101000";
        when "0111010010010" => rgb <= "101000";
        when "0111010010011" => rgb <= "101000";
        when "0111010010100" => rgb <= "101000";
        when "0111010010101" => rgb <= "101000";
        when "0111010010110" => rgb <= "101000";
        when "0111010010111" => rgb <= "101000";
        when "0111010011000" => rgb <= "101000";
        when "0111010011001" => rgb <= "101000";
        when "0111010011010" => rgb <= "101000";
        when "0111010011011" => rgb <= "000000";
        when "0111010011100" => rgb <= "100110";
        when "0111010011101" => rgb <= "100110";
        when "0111010011110" => rgb <= "100110";
        when "0111010011111" => rgb <= "100110";
        when "0111010100000" => rgb <= "000000";
        when "0111010100101" => rgb <= "000000";
        when "0111010100110" => rgb <= "100110";
        when "0111010100111" => rgb <= "100110";
        when "0111010101000" => rgb <= "100110";
        when "0111010101001" => rgb <= "100110";
        when "0111010101010" => rgb <= "000000";
        when "0111010101011" => rgb <= "100000";
        when "0111010101100" => rgb <= "100000";
        when "0111010101101" => rgb <= "100000";
        when "0111010101110" => rgb <= "100000";
        when "0111010101111" => rgb <= "100000";
        when "0111010110000" => rgb <= "100000";
        when "0111010110001" => rgb <= "100000";
        when "0111010110010" => rgb <= "100000";
        when "0111010110011" => rgb <= "100000";
        when "0111010110100" => rgb <= "100000";
        when "0111010110101" => rgb <= "000000";
        when "0111010110110" => rgb <= "101000";
        when "0111010110111" => rgb <= "101000";
        when "0111010111000" => rgb <= "101000";
        when "0111010111001" => rgb <= "101000";
        when "0111010111010" => rgb <= "101000";
        when "0111010111011" => rgb <= "101000";
        when "0111010111100" => rgb <= "101000";
        when "0111010111101" => rgb <= "101000";
        when "0111010111110" => rgb <= "101000";
        when "0111010111111" => rgb <= "101000";
        when "0111011000000" => rgb <= "000000";
        when "0111011000001" => rgb <= "000000";
        when "0111100001110" => rgb <= "000000";
        when "0111100001111" => rgb <= "000000";
        when "0111100010000" => rgb <= "101000";
        when "0111100010001" => rgb <= "101000";
        when "0111100010010" => rgb <= "101000";
        when "0111100010011" => rgb <= "101000";
        when "0111100010100" => rgb <= "101000";
        when "0111100010101" => rgb <= "101000";
        when "0111100010110" => rgb <= "101000";
        when "0111100010111" => rgb <= "101000";
        when "0111100011000" => rgb <= "101000";
        when "0111100011001" => rgb <= "101000";
        when "0111100011010" => rgb <= "101000";
        when "0111100011011" => rgb <= "000000";
        when "0111100011100" => rgb <= "100110";
        when "0111100011101" => rgb <= "100110";
        when "0111100011110" => rgb <= "100110";
        when "0111100011111" => rgb <= "100110";
        when "0111100100000" => rgb <= "100110";
        when "0111100100001" => rgb <= "000000";
        when "0111100100101" => rgb <= "000000";
        when "0111100100110" => rgb <= "100110";
        when "0111100100111" => rgb <= "100110";
        when "0111100101000" => rgb <= "100110";
        when "0111100101001" => rgb <= "100110";
        when "0111100101010" => rgb <= "000000";
        when "0111100101011" => rgb <= "100000";
        when "0111100101100" => rgb <= "100000";
        when "0111100101101" => rgb <= "100000";
        when "0111100101110" => rgb <= "100000";
        when "0111100101111" => rgb <= "100000";
        when "0111100110000" => rgb <= "100000";
        when "0111100110001" => rgb <= "100000";
        when "0111100110010" => rgb <= "100000";
        when "0111100110011" => rgb <= "100000";
        when "0111100110100" => rgb <= "100000";
        when "0111100110101" => rgb <= "000000";
        when "0111100110110" => rgb <= "101000";
        when "0111100110111" => rgb <= "101000";
        when "0111100111000" => rgb <= "101000";
        when "0111100111001" => rgb <= "101000";
        when "0111100111010" => rgb <= "000000";
        when "0111100111011" => rgb <= "000000";
        when "0111100111100" => rgb <= "000000";
        when "0111100111101" => rgb <= "101000";
        when "0111100111110" => rgb <= "101000";
        when "0111100111111" => rgb <= "101000";
        when "0111101000000" => rgb <= "101000";
        when "0111101000001" => rgb <= "000000";
        when "0111110001111" => rgb <= "000000";
        when "0111110010000" => rgb <= "000000";
        when "0111110010001" => rgb <= "101000";
        when "0111110010010" => rgb <= "101000";
        when "0111110010011" => rgb <= "101000";
        when "0111110010100" => rgb <= "101000";
        when "0111110010101" => rgb <= "101000";
        when "0111110010110" => rgb <= "101000";
        when "0111110010111" => rgb <= "101000";
        when "0111110011000" => rgb <= "101000";
        when "0111110011001" => rgb <= "101000";
        when "0111110011010" => rgb <= "101000";
        when "0111110011011" => rgb <= "000000";
        when "0111110011100" => rgb <= "100110";
        when "0111110011101" => rgb <= "100110";
        when "0111110011110" => rgb <= "100110";
        when "0111110011111" => rgb <= "100110";
        when "0111110100000" => rgb <= "100110";
        when "0111110100001" => rgb <= "000000";
        when "0111110100101" => rgb <= "000000";
        when "0111110100110" => rgb <= "100110";
        when "0111110100111" => rgb <= "100110";
        when "0111110101000" => rgb <= "100110";
        when "0111110101001" => rgb <= "100110";
        when "0111110101010" => rgb <= "000000";
        when "0111110101011" => rgb <= "100000";
        when "0111110101100" => rgb <= "100000";
        when "0111110101101" => rgb <= "100000";
        when "0111110101110" => rgb <= "100000";
        when "0111110101111" => rgb <= "100000";
        when "0111110110000" => rgb <= "100000";
        when "0111110110001" => rgb <= "100000";
        when "0111110110010" => rgb <= "000000";
        when "0111110110011" => rgb <= "000000";
        when "0111110110100" => rgb <= "000000";
        when "0111110110101" => rgb <= "000000";
        when "0111110110110" => rgb <= "101000";
        when "0111110110111" => rgb <= "101000";
        when "0111110111000" => rgb <= "101000";
        when "0111110111001" => rgb <= "000000";
        when "0111110111100" => rgb <= "000000";
        when "0111110111101" => rgb <= "101000";
        when "0111110111110" => rgb <= "101000";
        when "0111110111111" => rgb <= "101000";
        when "0111111000000" => rgb <= "101000";
        when "0111111000001" => rgb <= "000000";
        when "1000000010001" => rgb <= "000000";
        when "1000000010010" => rgb <= "101000";
        when "1000000010011" => rgb <= "101000";
        when "1000000010100" => rgb <= "101000";
        when "1000000010101" => rgb <= "101000";
        when "1000000010110" => rgb <= "101000";
        when "1000000010111" => rgb <= "101000";
        when "1000000011000" => rgb <= "101000";
        when "1000000011001" => rgb <= "101000";
        when "1000000011010" => rgb <= "101000";
        when "1000000011011" => rgb <= "101000";
        when "1000000011100" => rgb <= "000000";
        when "1000000011101" => rgb <= "100110";
        when "1000000011110" => rgb <= "100110";
        when "1000000011111" => rgb <= "100110";
        when "1000000100000" => rgb <= "100110";
        when "1000000100001" => rgb <= "000000";
        when "1000000100100" => rgb <= "000000";
        when "1000000100101" => rgb <= "100110";
        when "1000000100110" => rgb <= "100110";
        when "1000000100111" => rgb <= "100110";
        when "1000000101000" => rgb <= "100110";
        when "1000000101001" => rgb <= "100110";
        when "1000000101010" => rgb <= "000000";
        when "1000000101011" => rgb <= "100000";
        when "1000000101100" => rgb <= "100000";
        when "1000000101101" => rgb <= "100000";
        when "1000000101110" => rgb <= "000000";
        when "1000000101111" => rgb <= "000000";
        when "1000000110000" => rgb <= "000000";
        when "1000000110001" => rgb <= "000000";
        when "1000000110101" => rgb <= "000000";
        when "1000000110110" => rgb <= "101000";
        when "1000000110111" => rgb <= "101000";
        when "1000000111000" => rgb <= "101000";
        when "1000000111001" => rgb <= "101000";
        when "1000000111010" => rgb <= "000000";
        when "1000000111011" => rgb <= "000000";
        when "1000000111100" => rgb <= "000000";
        when "1000000111101" => rgb <= "101000";
        when "1000000111110" => rgb <= "101000";
        when "1000000111111" => rgb <= "101000";
        when "1000001000000" => rgb <= "101000";
        when "1000001000001" => rgb <= "000000";
        when "1000010010010" => rgb <= "000000";
        when "1000010010011" => rgb <= "000000";
        when "1000010010100" => rgb <= "101000";
        when "1000010010101" => rgb <= "101000";
        when "1000010010110" => rgb <= "101000";
        when "1000010010111" => rgb <= "101000";
        when "1000010011000" => rgb <= "101000";
        when "1000010011001" => rgb <= "101000";
        when "1000010011010" => rgb <= "101000";
        when "1000010011011" => rgb <= "101000";
        when "1000010011100" => rgb <= "000000";
        when "1000010011101" => rgb <= "000000";
        when "1000010011110" => rgb <= "100110";
        when "1000010011111" => rgb <= "100110";
        when "1000010100000" => rgb <= "100110";
        when "1000010100001" => rgb <= "000000";
        when "1000010100100" => rgb <= "000000";
        when "1000010100101" => rgb <= "100110";
        when "1000010100110" => rgb <= "100110";
        when "1000010100111" => rgb <= "100110";
        when "1000010101000" => rgb <= "100110";
        when "1000010101001" => rgb <= "000000";
        when "1000010101010" => rgb <= "100000";
        when "1000010101011" => rgb <= "100000";
        when "1000010101100" => rgb <= "100000";
        when "1000010101101" => rgb <= "000000";
        when "1000010110101" => rgb <= "000000";
        when "1000010110110" => rgb <= "101000";
        when "1000010110111" => rgb <= "101000";
        when "1000010111000" => rgb <= "101000";
        when "1000010111001" => rgb <= "101000";
        when "1000010111010" => rgb <= "101000";
        when "1000010111011" => rgb <= "101000";
        when "1000010111100" => rgb <= "101000";
        when "1000010111101" => rgb <= "101000";
        when "1000010111110" => rgb <= "101000";
        when "1000010111111" => rgb <= "101000";
        when "1000011000000" => rgb <= "101000";
        when "1000011000001" => rgb <= "000000";
        when "1000100010011" => rgb <= "000000";
        when "1000100010100" => rgb <= "000000";
        when "1000100010101" => rgb <= "101000";
        when "1000100010110" => rgb <= "101000";
        when "1000100010111" => rgb <= "101000";
        when "1000100011000" => rgb <= "101000";
        when "1000100011001" => rgb <= "101000";
        when "1000100011010" => rgb <= "101000";
        when "1000100011011" => rgb <= "101000";
        when "1000100011100" => rgb <= "101000";
        when "1000100011101" => rgb <= "000000";
        when "1000100011110" => rgb <= "100110";
        when "1000100011111" => rgb <= "100110";
        when "1000100100000" => rgb <= "100110";
        when "1000100100001" => rgb <= "100110";
        when "1000100100010" => rgb <= "000000";
        when "1000100100100" => rgb <= "000000";
        when "1000100100101" => rgb <= "100110";
        when "1000100100110" => rgb <= "100110";
        when "1000100100111" => rgb <= "100110";
        when "1000100101000" => rgb <= "100110";
        when "1000100101001" => rgb <= "000000";
        when "1000100101010" => rgb <= "100000";
        when "1000100101011" => rgb <= "100000";
        when "1000100101100" => rgb <= "100000";
        when "1000100101101" => rgb <= "100000";
        when "1000100101110" => rgb <= "000000";
        when "1000100101111" => rgb <= "000000";
        when "1000100110000" => rgb <= "000000";
        when "1000100110101" => rgb <= "000000";
        when "1000100110110" => rgb <= "101000";
        when "1000100110111" => rgb <= "101000";
        when "1000100111000" => rgb <= "101000";
        when "1000100111001" => rgb <= "101000";
        when "1000100111010" => rgb <= "101000";
        when "1000100111011" => rgb <= "101000";
        when "1000100111100" => rgb <= "101000";
        when "1000100111101" => rgb <= "101000";
        when "1000100111110" => rgb <= "101000";
        when "1000100111111" => rgb <= "101000";
        when "1000101000000" => rgb <= "000000";
        when "1000110010101" => rgb <= "000000";
        when "1000110010110" => rgb <= "101000";
        when "1000110010111" => rgb <= "101000";
        when "1000110011000" => rgb <= "101000";
        when "1000110011001" => rgb <= "101000";
        when "1000110011010" => rgb <= "101000";
        when "1000110011011" => rgb <= "101000";
        when "1000110011100" => rgb <= "101000";
        when "1000110011101" => rgb <= "000000";
        when "1000110011110" => rgb <= "100110";
        when "1000110011111" => rgb <= "100110";
        when "1000110100000" => rgb <= "100110";
        when "1000110100001" => rgb <= "100110";
        when "1000110100010" => rgb <= "000000";
        when "1000110100011" => rgb <= "000000";
        when "1000110100100" => rgb <= "100110";
        when "1000110100101" => rgb <= "100110";
        when "1000110100110" => rgb <= "100110";
        when "1000110100111" => rgb <= "100110";
        when "1000110101000" => rgb <= "100110";
        when "1000110101001" => rgb <= "000000";
        when "1000110101010" => rgb <= "100000";
        when "1000110101011" => rgb <= "100000";
        when "1000110101100" => rgb <= "100000";
        when "1000110101101" => rgb <= "100000";
        when "1000110101110" => rgb <= "100000";
        when "1000110101111" => rgb <= "100000";
        when "1000110110000" => rgb <= "100000";
        when "1000110110001" => rgb <= "000000";
        when "1000110110101" => rgb <= "000000";
        when "1000110110110" => rgb <= "101000";
        when "1000110110111" => rgb <= "101000";
        when "1000110111000" => rgb <= "101000";
        when "1000110111001" => rgb <= "101000";
        when "1000110111010" => rgb <= "101000";
        when "1000110111011" => rgb <= "101000";
        when "1000110111100" => rgb <= "101000";
        when "1000110111101" => rgb <= "101000";
        when "1000110111110" => rgb <= "101000";
        when "1000110111111" => rgb <= "101000";
        when "1000111000000" => rgb <= "000000";
        when "1000111000001" => rgb <= "000000";
        when "1001000010101" => rgb <= "000000";
        when "1001000010110" => rgb <= "101000";
        when "1001000010111" => rgb <= "101000";
        when "1001000011000" => rgb <= "101000";
        when "1001000011001" => rgb <= "101000";
        when "1001000011010" => rgb <= "101000";
        when "1001000011011" => rgb <= "101000";
        when "1001000011100" => rgb <= "101000";
        when "1001000011101" => rgb <= "000000";
        when "1001000011110" => rgb <= "100110";
        when "1001000011111" => rgb <= "100110";
        when "1001000100000" => rgb <= "100110";
        when "1001000100001" => rgb <= "100110";
        when "1001000100010" => rgb <= "100110";
        when "1001000100011" => rgb <= "100110";
        when "1001000100100" => rgb <= "100110";
        when "1001000100101" => rgb <= "100110";
        when "1001000100110" => rgb <= "100110";
        when "1001000100111" => rgb <= "100110";
        when "1001000101000" => rgb <= "000000";
        when "1001000101001" => rgb <= "000000";
        when "1001000101010" => rgb <= "100000";
        when "1001000101011" => rgb <= "100000";
        when "1001000101100" => rgb <= "100000";
        when "1001000101101" => rgb <= "100000";
        when "1001000101110" => rgb <= "100000";
        when "1001000101111" => rgb <= "100000";
        when "1001000110000" => rgb <= "100000";
        when "1001000110001" => rgb <= "000000";
        when "1001000110101" => rgb <= "000000";
        when "1001000110110" => rgb <= "101000";
        when "1001000110111" => rgb <= "101000";
        when "1001000111000" => rgb <= "101000";
        when "1001000111001" => rgb <= "101000";
        when "1001000111010" => rgb <= "000000";
        when "1001000111011" => rgb <= "000000";
        when "1001000111100" => rgb <= "000000";
        when "1001000111101" => rgb <= "000000";
        when "1001000111110" => rgb <= "101000";
        when "1001000111111" => rgb <= "101000";
        when "1001001000000" => rgb <= "101000";
        when "1001001000001" => rgb <= "000000";
        when "1001010010100" => rgb <= "000000";
        when "1001010010101" => rgb <= "101000";
        when "1001010010110" => rgb <= "101000";
        when "1001010010111" => rgb <= "101000";
        when "1001010011000" => rgb <= "101000";
        when "1001010011001" => rgb <= "101000";
        when "1001010011010" => rgb <= "101000";
        when "1001010011011" => rgb <= "101000";
        when "1001010011100" => rgb <= "101000";
        when "1001010011101" => rgb <= "000000";
        when "1001010011110" => rgb <= "100110";
        when "1001010011111" => rgb <= "100110";
        when "1001010100000" => rgb <= "100110";
        when "1001010100001" => rgb <= "100110";
        when "1001010100010" => rgb <= "100110";
        when "1001010100011" => rgb <= "100110";
        when "1001010100100" => rgb <= "100110";
        when "1001010100101" => rgb <= "100110";
        when "1001010100110" => rgb <= "100110";
        when "1001010100111" => rgb <= "100110";
        when "1001010101000" => rgb <= "000000";
        when "1001010101001" => rgb <= "000000";
        when "1001010101010" => rgb <= "100000";
        when "1001010101011" => rgb <= "100000";
        when "1001010101100" => rgb <= "100000";
        when "1001010101101" => rgb <= "100000";
        when "1001010101110" => rgb <= "000000";
        when "1001010101111" => rgb <= "000000";
        when "1001010110000" => rgb <= "000000";
        when "1001010110001" => rgb <= "000000";
        when "1001010110101" => rgb <= "000000";
        when "1001010110110" => rgb <= "101000";
        when "1001010110111" => rgb <= "101000";
        when "1001010111000" => rgb <= "101000";
        when "1001010111001" => rgb <= "101000";
        when "1001010111010" => rgb <= "000000";
        when "1001010111110" => rgb <= "000000";
        when "1001010111111" => rgb <= "101000";
        when "1001011000000" => rgb <= "101000";
        when "1001011000001" => rgb <= "101000";
        when "1001011000010" => rgb <= "000000";
        when "1001100010011" => rgb <= "000000";
        when "1001100010100" => rgb <= "101000";
        when "1001100010101" => rgb <= "101000";
        when "1001100010110" => rgb <= "101000";
        when "1001100010111" => rgb <= "101000";
        when "1001100011000" => rgb <= "101000";
        when "1001100011001" => rgb <= "101000";
        when "1001100011010" => rgb <= "101000";
        when "1001100011011" => rgb <= "101000";
        when "1001100011100" => rgb <= "101000";
        when "1001100011101" => rgb <= "101000";
        when "1001100011110" => rgb <= "000000";
        when "1001100011111" => rgb <= "100110";
        when "1001100100000" => rgb <= "100110";
        when "1001100100001" => rgb <= "100110";
        when "1001100100010" => rgb <= "100110";
        when "1001100100011" => rgb <= "100110";
        when "1001100100100" => rgb <= "100110";
        when "1001100100101" => rgb <= "100110";
        when "1001100100110" => rgb <= "100110";
        when "1001100100111" => rgb <= "000000";
        when "1001100101001" => rgb <= "000000";
        when "1001100101010" => rgb <= "100000";
        when "1001100101011" => rgb <= "100000";
        when "1001100101100" => rgb <= "100000";
        when "1001100101101" => rgb <= "100000";
        when "1001100101110" => rgb <= "000000";
        when "1001100101111" => rgb <= "000000";
        when "1001100110101" => rgb <= "000000";
        when "1001100110110" => rgb <= "101000";
        when "1001100110111" => rgb <= "101000";
        when "1001100111000" => rgb <= "101000";
        when "1001100111001" => rgb <= "101000";
        when "1001100111010" => rgb <= "000000";
        when "1001100111110" => rgb <= "000000";
        when "1001100111111" => rgb <= "101000";
        when "1001101000000" => rgb <= "101000";
        when "1001101000001" => rgb <= "101000";
        when "1001101000010" => rgb <= "000000";
        when "1001101000011" => rgb <= "000000";
        when "1001110010010" => rgb <= "000000";
        when "1001110010011" => rgb <= "101000";
        when "1001110010100" => rgb <= "101000";
        when "1001110010101" => rgb <= "101000";
        when "1001110010110" => rgb <= "101000";
        when "1001110010111" => rgb <= "101000";
        when "1001110011000" => rgb <= "101000";
        when "1001110011001" => rgb <= "101000";
        when "1001110011010" => rgb <= "101000";
        when "1001110011011" => rgb <= "101000";
        when "1001110011100" => rgb <= "101000";
        when "1001110011101" => rgb <= "000000";
        when "1001110011110" => rgb <= "000000";
        when "1001110011111" => rgb <= "100110";
        when "1001110100000" => rgb <= "100110";
        when "1001110100001" => rgb <= "100110";
        when "1001110100010" => rgb <= "100110";
        when "1001110100011" => rgb <= "100110";
        when "1001110100100" => rgb <= "100110";
        when "1001110100101" => rgb <= "100110";
        when "1001110100110" => rgb <= "100110";
        when "1001110100111" => rgb <= "000000";
        when "1001110101001" => rgb <= "000000";
        when "1001110101010" => rgb <= "100000";
        when "1001110101011" => rgb <= "100000";
        when "1001110101100" => rgb <= "100000";
        when "1001110101101" => rgb <= "100000";
        when "1001110101110" => rgb <= "100000";
        when "1001110101111" => rgb <= "000000";
        when "1001110110000" => rgb <= "000000";
        when "1001110110001" => rgb <= "000000";
        when "1001110110010" => rgb <= "000000";
        when "1001110110011" => rgb <= "000000";
        when "1001110110100" => rgb <= "000000";
        when "1001110110101" => rgb <= "000000";
        when "1001110110110" => rgb <= "000000";
        when "1001110110111" => rgb <= "101000";
        when "1001110111000" => rgb <= "101000";
        when "1001110111001" => rgb <= "101000";
        when "1001110111010" => rgb <= "000000";
        when "1001110111110" => rgb <= "000000";
        when "1001110111111" => rgb <= "000000";
        when "1001111000000" => rgb <= "101000";
        when "1001111000001" => rgb <= "101000";
        when "1001111000010" => rgb <= "101000";
        when "1001111000011" => rgb <= "000000";
        when "1010000010001" => rgb <= "000000";
        when "1010000010010" => rgb <= "101000";
        when "1010000010011" => rgb <= "101000";
        when "1010000010100" => rgb <= "101000";
        when "1010000010101" => rgb <= "101000";
        when "1010000010110" => rgb <= "101000";
        when "1010000010111" => rgb <= "101000";
        when "1010000011000" => rgb <= "101000";
        when "1010000011001" => rgb <= "101000";
        when "1010000011010" => rgb <= "101000";
        when "1010000011011" => rgb <= "101000";
        when "1010000011100" => rgb <= "101000";
        when "1010000011101" => rgb <= "000000";
        when "1010000011111" => rgb <= "000000";
        when "1010000100000" => rgb <= "100110";
        when "1010000100001" => rgb <= "100110";
        when "1010000100010" => rgb <= "100110";
        when "1010000100011" => rgb <= "100110";
        when "1010000100100" => rgb <= "100110";
        when "1010000100101" => rgb <= "100110";
        when "1010000100110" => rgb <= "000000";
        when "1010000100111" => rgb <= "000000";
        when "1010000101010" => rgb <= "000000";
        when "1010000101011" => rgb <= "100000";
        when "1010000101100" => rgb <= "100000";
        when "1010000101101" => rgb <= "100000";
        when "1010000101110" => rgb <= "100000";
        when "1010000101111" => rgb <= "100000";
        when "1010000110000" => rgb <= "100000";
        when "1010000110001" => rgb <= "100000";
        when "1010000110010" => rgb <= "100000";
        when "1010000110011" => rgb <= "100000";
        when "1010000110100" => rgb <= "100000";
        when "1010000110101" => rgb <= "100000";
        when "1010000110110" => rgb <= "000000";
        when "1010000110111" => rgb <= "000000";
        when "1010000111000" => rgb <= "101000";
        when "1010000111001" => rgb <= "101000";
        when "1010000111010" => rgb <= "000000";
        when "1010000111111" => rgb <= "000000";
        when "1010001000000" => rgb <= "101000";
        when "1010001000001" => rgb <= "101000";
        when "1010001000010" => rgb <= "101000";
        when "1010001000011" => rgb <= "000000";
        when "1010010010000" => rgb <= "000000";
        when "1010010010001" => rgb <= "101000";
        when "1010010010010" => rgb <= "101000";
        when "1010010010011" => rgb <= "101000";
        when "1010010010100" => rgb <= "101000";
        when "1010010010101" => rgb <= "101000";
        when "1010010010110" => rgb <= "101000";
        when "1010010010111" => rgb <= "101000";
        when "1010010011000" => rgb <= "101000";
        when "1010010011001" => rgb <= "101000";
        when "1010010011010" => rgb <= "101000";
        when "1010010011011" => rgb <= "101000";
        when "1010010011100" => rgb <= "000000";
        when "1010010011111" => rgb <= "000000";
        when "1010010100000" => rgb <= "000000";
        when "1010010100001" => rgb <= "100110";
        when "1010010100010" => rgb <= "100110";
        when "1010010100011" => rgb <= "100110";
        when "1010010100100" => rgb <= "100110";
        when "1010010100101" => rgb <= "100110";
        when "1010010100110" => rgb <= "000000";
        when "1010010101010" => rgb <= "000000";
        when "1010010101011" => rgb <= "100000";
        when "1010010101100" => rgb <= "100000";
        when "1010010101101" => rgb <= "100000";
        when "1010010101110" => rgb <= "100000";
        when "1010010101111" => rgb <= "100000";
        when "1010010110000" => rgb <= "100000";
        when "1010010110001" => rgb <= "100000";
        when "1010010110010" => rgb <= "100000";
        when "1010010110011" => rgb <= "100000";
        when "1010010110100" => rgb <= "100000";
        when "1010010110101" => rgb <= "100000";
        when "1010010110110" => rgb <= "100000";
        when "1010010110111" => rgb <= "000000";
        when "1010010111000" => rgb <= "101000";
        when "1010010111001" => rgb <= "101000";
        when "1010010111010" => rgb <= "000000";
        when "1010010111111" => rgb <= "000000";
        when "1010011000000" => rgb <= "101000";
        when "1010011000001" => rgb <= "101000";
        when "1010011000010" => rgb <= "101000";
        when "1010011000011" => rgb <= "000000";
        when "1010100001110" => rgb <= "000000";
        when "1010100001111" => rgb <= "000000";
        when "1010100010000" => rgb <= "101000";
        when "1010100010001" => rgb <= "101000";
        when "1010100010010" => rgb <= "101000";
        when "1010100010011" => rgb <= "101000";
        when "1010100010100" => rgb <= "101000";
        when "1010100010101" => rgb <= "101000";
        when "1010100010110" => rgb <= "101000";
        when "1010100010111" => rgb <= "101000";
        when "1010100011000" => rgb <= "101000";
        when "1010100011001" => rgb <= "101000";
        when "1010100011010" => rgb <= "101000";
        when "1010100011011" => rgb <= "000000";
        when "1010100100000" => rgb <= "000000";
        when "1010100100001" => rgb <= "000000";
        when "1010100100010" => rgb <= "100110";
        when "1010100100011" => rgb <= "100110";
        when "1010100100100" => rgb <= "100110";
        when "1010100100101" => rgb <= "000000";
        when "1010100101010" => rgb <= "000000";
        when "1010100101011" => rgb <= "100000";
        when "1010100101100" => rgb <= "100000";
        when "1010100101101" => rgb <= "100000";
        when "1010100101110" => rgb <= "100000";
        when "1010100101111" => rgb <= "100000";
        when "1010100110000" => rgb <= "100000";
        when "1010100110001" => rgb <= "100000";
        when "1010100110010" => rgb <= "100000";
        when "1010100110011" => rgb <= "100000";
        when "1010100110100" => rgb <= "100000";
        when "1010100110101" => rgb <= "100000";
        when "1010100110110" => rgb <= "100000";
        when "1010100110111" => rgb <= "000000";
        when "1010100111000" => rgb <= "101000";
        when "1010100111001" => rgb <= "101000";
        when "1010100111010" => rgb <= "000000";
        when "1010100111111" => rgb <= "000000";
        when "1010101000000" => rgb <= "000000";
        when "1010101000001" => rgb <= "101000";
        when "1010101000010" => rgb <= "101000";
        when "1010101000011" => rgb <= "000000";
        when "1010110001111" => rgb <= "000000";
        when "1010110010000" => rgb <= "101000";
        when "1010110010001" => rgb <= "101000";
        when "1010110010010" => rgb <= "101000";
        when "1010110010011" => rgb <= "101000";
        when "1010110010100" => rgb <= "101000";
        when "1010110010101" => rgb <= "101000";
        when "1010110010110" => rgb <= "101000";
        when "1010110010111" => rgb <= "101000";
        when "1010110011000" => rgb <= "101000";
        when "1010110011001" => rgb <= "101000";
        when "1010110011010" => rgb <= "000000";
        when "1010110100001" => rgb <= "000000";
        when "1010110100010" => rgb <= "100110";
        when "1010110100011" => rgb <= "100110";
        when "1010110100100" => rgb <= "100110";
        when "1010110100101" => rgb <= "000000";
        when "1010110101010" => rgb <= "000000";
        when "1010110101011" => rgb <= "100000";
        when "1010110101100" => rgb <= "100000";
        when "1010110101101" => rgb <= "100000";
        when "1010110101110" => rgb <= "100000";
        when "1010110101111" => rgb <= "100000";
        when "1010110110000" => rgb <= "100000";
        when "1010110110001" => rgb <= "100000";
        when "1010110110010" => rgb <= "100000";
        when "1010110110011" => rgb <= "100000";
        when "1010110110100" => rgb <= "100000";
        when "1010110110101" => rgb <= "000000";
        when "1010110110110" => rgb <= "000000";
        when "1010110110111" => rgb <= "000000";
        when "1010110111000" => rgb <= "101000";
        when "1010110111001" => rgb <= "000000";
        when "1010110111010" => rgb <= "000000";
        when "1010111000000" => rgb <= "000000";
        when "1010111000001" => rgb <= "101000";
        when "1010111000010" => rgb <= "000000";
        when "1010111000011" => rgb <= "000000";
        when "1011000010000" => rgb <= "000000";
        when "1011000010001" => rgb <= "000000";
        when "1011000010010" => rgb <= "101000";
        when "1011000010011" => rgb <= "101000";
        when "1011000010100" => rgb <= "101000";
        when "1011000010101" => rgb <= "101000";
        when "1011000010110" => rgb <= "101000";
        when "1011000010111" => rgb <= "000000";
        when "1011000011000" => rgb <= "000000";
        when "1011000011001" => rgb <= "000000";
        when "1011000100010" => rgb <= "000000";
        when "1011000100011" => rgb <= "000000";
        when "1011000100100" => rgb <= "000000";
        when "1011000100101" => rgb <= "000000";
        when "1011000101011" => rgb <= "000000";
        when "1011000101100" => rgb <= "000000";
        when "1011000101101" => rgb <= "000000";
        when "1011000101110" => rgb <= "000000";
        when "1011000101111" => rgb <= "000000";
        when "1011000110000" => rgb <= "000000";
        when "1011000110001" => rgb <= "000000";
        when "1011000110010" => rgb <= "000000";
        when "1011000110011" => rgb <= "000000";
        when "1011000110100" => rgb <= "000000";
        when "1011000110101" => rgb <= "000000";
        when "1011000110111" => rgb <= "000000";
        when "1011000111000" => rgb <= "000000";
        when "1011000111001" => rgb <= "000000";
        when "1011001000001" => rgb <= "000000";
        when "1011001000010" => rgb <= "000000";
        when "1011010010010" => rgb <= "000000";
        when "1011010010011" => rgb <= "000000";
        when "1011010010100" => rgb <= "000000";
        when "1011010010101" => rgb <= "000000";
        when "1011010010110" => rgb <= "000000";
        when others => rgb <= "001000";
            end case;
   end process;
end Behavioral;

